`timescale 1ns/1ps

module adder_32_tb;

  // Parameters
  localparam WIDTH = 32;

  // Signals
  reg [WIDTH-1:0] a;
  reg [WIDTH-1:0] b;
  wire [WIDTH-1:0] y;

  // Instantiate the adder_32 module
  adder_32 #(WIDTH) dut (
    .a(a),
    .b(b),
    .y(y)
  );

  // Test cases
  initial begin
    // Test 1: Add two positive numbers
    a = 32'h12345678;
    b = 32'h87654321;
    #10;
    $display("Test 1: Add two positive numbers");
    $display("a: %h", a);
    $display("b: %h", b);
    $display("y (a + b): %h", y);

    // Test 2: Add a positive and a negative number
    a = 32'h12345678;
    b = 32'h87654321; // Negative number
    #10;
    $display("Test 2: Add a positive and a negative number");
    $display("a: %h", a);
    $display("b: %h", b);
    $display("y (a + b): %h", y);

    // Test 3: Add two negative numbers
    a = 32'h12345678; // Negative number
    b = 32'h87654321; // Negative number
    #10;
    $display("Test 3: Add two negative numbers");
    $display("a: %h", a);
    $display("b: %h", b);
    $display("y (a + b): %h", y);

    // Add more test cases...

    // Finish the simulation
    $finish;
  end

endmodule

`timescale 1ns/1ps

module RegFiles_tb;

  // Parameters
  localparam DATA_WIDTH = 32;
  localparam ADDRESS_WIDTH = 5;
  localparam NUM_REGS = 32;

  // Signals
  reg clk = 0;
  reg rst = 0;
  reg RegWrite = 0;
  reg [ADDRESS_WIDTH-1:0] rg_wrt_dest;
  reg [ADDRESS_WIDTH-1:0] rs1;
  reg [ADDRESS_WIDTH-1:0] rs2;
  reg [DATA_WIDTH-1:0] rg_wrt_data;
  wire [DATA_WIDTH-1:0] read_reg1;
  wire [DATA_WIDTH-1:0] read_reg2;

  // Instantiate the RegFiles module
  RegFiles #(DATA_WIDTH, ADDRESS_WIDTH, NUM_REGS) dut (
    .clk(clk),
    .rst(rst),
    .RegWrite(RegWrite),
    .rg_wrt_dest(rg_wrt_dest),
    .rs1(rs1),
    .rs2(rs2),
    .rg_wrt_data(rg_wrt_data),
    .read_reg1(read_reg1),
    .read_reg2(read_reg2)
  );

  // Clock generation
  always begin
    #5 clk = ~clk;
  end

  // Test cases
  initial begin
    // Test 1: Write to and read from a register
    rst = 1'b0;
    RegWrite = 1'b1;
    rg_wrt_dest = 5'b00100; // Write to register 4
    rg_wrt_data = 32'h12345678; // Data to write
    rs1 = 5'b00001; // Read from register 1
    rs2 = 5'b00100; // Read from register 4
	 
    #10;
    $display("Test 1: Write to and read from a register");
    $display("Write Data: %h", rg_wrt_data);
    $display("Read Register 1: %h", read_reg1);
    $display("Read Register 2: %h", read_reg2);

    // Add more test cases...

    // Finish the simulation
    $finish;
  end

endmodule
